// Module: Program Counter
// Author: M.M.C.J.Bandara - 180065C
// xx/01/2022

module name(   
    input clk,                  // Clock

);

always @ (posedge clk)
begin

end

endmodule